/* Advanced Digital Design 2025

Title: shiftreg.v 
Description: This HDL code is an example of basics
definitions of modules which involves I/O. 
Author: Corvalan, Abel.

*/

module shiftreg(
    output [] outshif,
    input  [] 
);

endmodule