/* Advanced Digital Design 2025

Title: shiftreg.v 
Description: This HDL code is an example of basics
definitions of modules which involves I/O. 
Author: Corvalan, Abel.

*/

module shiftreg(
    output [3:0] o_led,

    input      i_valid, 
    input      i_reset,
    input        clock;
);

endmodule