/* Advanced Digital Design 2025

Title: count.v 
Description: This HDL code is an example of basics
definitions of modules which involves I/O. 
Author: Corvalan, Abel.

*/

module count (
    output      o_valid,
    
    input [2:0] i_sw   ,
    input       i_reset,
    input       clock  
);

endmodule